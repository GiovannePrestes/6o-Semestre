library verilog;
use verilog.vl_types.all;
entity mem_4x16_vlg_vec_tst is
end mem_4x16_vlg_vec_tst;
