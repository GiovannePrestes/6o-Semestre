library verilog;
use verilog.vl_types.all;
entity Reg4bits_vlg_vec_tst is
end Reg4bits_vlg_vec_tst;
