library verilog;
use verilog.vl_types.all;
entity mem_4x16_vlg_check_tst is
    port(
        OUT_0           : in     vl_logic;
        OUT_1           : in     vl_logic;
        OUT_2           : in     vl_logic;
        OUT_3           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mem_4x16_vlg_check_tst;
