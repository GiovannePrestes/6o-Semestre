library verilog;
use verilog.vl_types.all;
entity bitBuffer_vlg_vec_tst is
end bitBuffer_vlg_vec_tst;
